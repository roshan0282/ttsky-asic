//`timescale 1ns / 1ps


// input 0-89 degree, Q0.8 [0,1] 0.004
//  - case: 90 = 256, handle outside this module
//  - dont forget to convert Q0.8 to Q8.8

// const fix sinTable[] = {
// 0,4,8,13,17,22,26,31,35,40,44,48,53,57,61,66,70,74,79,83,87,91,95,100,104,108,112,
// 116,120,124,128,131,135,139,143,146,150,154,157,161,164,167,171,174,177,181,184,187,
// 190,193,196,198,201,204,207,209,212,214,217,219,221,223,226,228,230,232,233,235,237,
// 238,240,242,243,244,246,247,248,249,250,251,252,252,253,254,254,255,255,255,255,255};



module sine_rom (
    input wire [6:0]  angle,
    output wire [7:0] value
);

  reg [7:0] mem;
  assign value = mem;

  always @(*) begin
    case(angle)
      0: mem = 0;
      1: mem = 4;
      2: mem = 8;
      3: mem = 13;
      4: mem = 17;
      5: mem = 22;
      6: mem = 26;
      7: mem = 31;
      8: mem = 35;
      9: mem = 40;
      10: mem = 44;
      11: mem = 48;
      12: mem = 53;
      13: mem = 57;
      14: mem = 61;
      15: mem = 66;
      16: mem = 70;
      17: mem = 74;
      18: mem = 79;
      19: mem = 83;
      20: mem = 87;
      21: mem = 91;
      22: mem = 95;
      23: mem = 100;
      24: mem = 104;
      25: mem = 108;
      26: mem = 112;
      27: mem = 116;
      28: mem = 120;
      29: mem = 124;
      30: mem = 128;
      31: mem = 131;
      32: mem = 135;
      33: mem = 139;
      34: mem = 143;
      35: mem = 146;
      36: mem = 150;
      37: mem = 154;
      38: mem = 157;
      39: mem = 161;
      40: mem = 164;
      41: mem = 167;
      42: mem = 171;
      43: mem = 174;
      44: mem = 177;
      45: mem = 181;
      46: mem = 184;
      47: mem = 187;
      48: mem = 190;
      49: mem = 193;
      50: mem = 196;
      51: mem = 198;
      52: mem = 201;
      53: mem = 204;
      54: mem = 207;
      55: mem = 209;
      56: mem = 212;
      57: mem = 214;
      58: mem = 217;
      59: mem = 219;
      60: mem = 221;
      61: mem = 223;
      62: mem = 226;
      63: mem = 228;
      64: mem = 230;
      65: mem = 232;
      66: mem = 233;
      67: mem = 235;
      68: mem = 237;
      69: mem = 238;
      70: mem = 240;
      71: mem = 242;
      72: mem = 243;
      73: mem = 244;
      74: mem = 246;
      75: mem = 247;
      76: mem = 248;
      77: mem = 249;
      78: mem = 250;
      79: mem = 251;
      80: mem = 252;
      81: mem = 252;
      82: mem = 253;
      83: mem = 254;
      84: mem = 254;
      85: mem = 255;
      86: mem = 255;
      87: mem = 255;
      88: mem = 255;
      89: mem = 255;
      default: mem = 0;
    endcase
  end




endmodule
